`timescale 1ns / 1ps
module opt_check2 (input a , input b , output y);
	assign y = a?1:b;
endmodule
